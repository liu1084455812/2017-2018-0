library verilog;
use verilog.vl_types.all;
entity PC is
    port(
        rst             : in     vl_logic;
        clk             : in     vl_logic;
        PCWrite         : in     vl_logic;
        nPC             : in     vl_logic_vector(31 downto 0);
        PC              : out    vl_logic_vector(31 downto 0)
    );
end PC;
